/*
 * Copyright 2018 Akifumi Fujita
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

import BasicTypes::*;
import RvTypes::*;
import Rv32Types::*;

import CacheTypes::*;

interface FetchAddrTranslateStageIF;
    logic valid;
    logic tlbFault;
    logic tlbMiss;
    vaddr_t pc_vaddr;
    paddr_t pc_paddr;

    modport ThisStage(
    output
        valid,
        tlbFault,
        tlbMiss,
        pc_vaddr,
        pc_paddr
    );

    modport NextStage(
    input
        valid,
        tlbFault,
        tlbMiss,
        pc_vaddr,
        pc_paddr
    );
endinterface
