/*
 * Copyright 2018 Akifumi Fujita
 * 
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 * 
 *     http://www.apache.org/licenses/LICENSE-2.0
 * 
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

import BasicTypes::*;
import RvTypes::*;
import Rv32Types::*;

import ProcessorTypes::*;

module BypassLogic(
    BypassLogicIF.BypassLogic bus,
    PipelineControllerIF.BypassLogic ctrl,
    input clk,
    input rst
);
    typedef logic [$clog2(BypassDepth)-1:0] _index_t;

    typedef struct packed {
        logic valid;
        reg_addr_t addr;
        word_t value;
    } PipelineEntry;

    // Functions
    function automatic _index_t encodeIndex(logic [BypassDepth-1:0] depth);
        for (int i = 0; i < BypassDepth; i++) begin
            if (depth[i]) begin
                return i;
            end
        end
        return 0;
    endfunction

    // Registers
    PipelineEntry pipeline[BypassDepth];

    // Wires
    logic loadHit[BypassReadPortCount];
    logic [BypassDepth-1:0] camHits[BypassReadPortCount];
    _index_t camIndex[BypassReadPortCount];

    // Bypass CAM
    always_comb begin
        for (int i = 0; i < BypassReadPortCount; i++) begin
            loadHit[i] = bus.loadWriteEnable && bus.loadWriteAddr == bus.readAddr[i];

            for (int j = 0; j < BypassDepth; j++) begin
                camHits[i][j] = pipeline[j].valid && (pipeline[j].addr == bus.readAddr[i]);
            end
            camIndex[i] = encodeIndex(camHits[i]);

            bus.hit[i] = |(camHits[i]) || loadHit[i];
            if (bus.readAddr[i] == '0) begin
                // zero register
                bus.readValue[i] = '0;
            end
            else if (loadHit[i]) begin
                bus.readValue[i] = bus.loadWriteValue;
            end
            else if (|(camHits[i])) begin
                bus.readValue[i] = pipeline[camIndex[i]].value;
            end
            else begin
                // bypass failure
                bus.readValue[i] = '0;
            end
        end
    end

    // Bypass Pipeline
    always_ff @(posedge clk) begin
        if (rst || ctrl.flush) begin
            for (int i = 0; i < BypassDepth; i++) begin
                pipeline[i] <= '0;
            end
        end
        else if (ctrl.stall) begin
            for (int i = 0; i < BypassDepth; i++) begin
                pipeline[i] <= pipeline[i];
            end
        end
        else begin
            pipeline[0].valid <= bus.writeEnable;
            pipeline[0].addr <= bus.writeAddr;
            pipeline[0].value <= bus.writeValue;
            
            if (bus.loadWriteEnable) begin
                pipeline[1].valid <= bus.loadWriteEnable;
                pipeline[1].addr <= bus.loadWriteAddr;
                pipeline[1].value <= bus.loadWriteValue;
            end
            else begin
                pipeline[1] <= pipeline[0];
            end
            
            for (int i = 2; i < BypassDepth; i++) begin
                pipeline[i] <= pipeline[i-1];
            end
        end
    end
endmodule
